
module moduleName (
    ports
);
    
endmodule