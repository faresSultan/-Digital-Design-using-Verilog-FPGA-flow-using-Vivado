module Q1_tb ();
    

    
endmodule