module moduleName (
    ports
);
    
endmodule
